library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity OutputIEEE_8_23_to_8_23 is
    port ( X : in  std_logic_vector(8+23+2 downto 0);
           R : out  std_logic_vector(31 downto 0)   );
end entity;

architecture arch of OutputIEEE_8_23_to_8_23 is
signal expX :  std_logic_vector(7 downto 0);
signal fracX :  std_logic_vector(22 downto 0);
signal exnX :  std_logic_vector(1 downto 0);
signal sX :  std_logic;
signal expZero :  std_logic;
signal sfracX :  std_logic_vector(22 downto 0);
signal fracR :  std_logic_vector(22 downto 0);
signal expR :  std_logic_vector(7 downto 0);
begin
    expX  <= X(30 downto 23);
    fracX  <= X(22 downto 0);
    exnX  <= X(33 downto 32);
    sX  <= X(31) when (exnX = "01" or exnX = "10" or exnX = "00") else '0';
    expZero  <= '1' when expX = (7 downto 0 => '0') else '0';
    -- since we have one more exponent value than IEEE (field 0...0, value emin-1),
    -- we can represent subnormal numbers whose mantissa field begins with a 1
    sfracX <= 
      (22 downto 0 => '0') when (exnX = "00") else
      '1' & fracX(22 downto 1) when (expZero = '1' and exnX = "01") else
      fracX when (exnX = "01") else 
      (22 downto 1 => '0') & exnX(0);
    fracR <= sfracX;
    expR <=  
      (7 downto 0 => '0') when (exnX = "00") else
      expX when (exnX = "01") else 
      (7 downto 0 => '1');
    R <= sX & expR & fracR; 
end architecture;